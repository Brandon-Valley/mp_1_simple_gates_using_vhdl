og_code_str,code,adv_value,real_value
6006491646202759848              
6006491646202730435              
6006491646202685902              
6006491646202707078              
6006491646204098450              
