
library ieee;
use ieee.std_logic_1164.all;


entity and_gate is
  port ( A: in std_logic;
         B: in std_logic;
         F: out std_logic);
end and_gate;

architecture behavior of and_gate is
  begin
    F <= A and B;
end behavior;

